module some_project;
    import some_published_dependency::*;
endmodule
