class some_class;

    function void do_some_other_thing();
      $display("doing some other thing");
    endfunction

endclass
