package some_published_dependency;
endpackage
