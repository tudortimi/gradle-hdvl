package dummy0;
  import dummy1::*;
endpackage
