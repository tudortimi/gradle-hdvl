package some_project;
endpackage
