package some_published_dependency;
    `include "some_class.svh"
    import "DPI-C" function void some_dpi_func();
endpackage
