package proj0;
endpackage
