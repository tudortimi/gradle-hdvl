package dummy1;
endpackage
