package tb;
endpackage
