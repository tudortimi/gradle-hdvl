package dummy2;
  import dummy1::*;
endpackage
