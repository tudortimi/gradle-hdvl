class some_class;

  function void do_some_thing();
    $display("doing some thing");
  endfunction

endclass
