class some_class;

    function bit is_working();
        return 1;
    endfunction

endclass
