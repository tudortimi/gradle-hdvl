package dummy0;
  import dummy1::*;
  import dummy2::*;
endpackage
