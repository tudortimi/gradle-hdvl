package utils0;
endpackage
