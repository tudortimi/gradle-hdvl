package utils;
endpackage
