package some_package;
endpackage
