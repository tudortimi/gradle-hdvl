package test_utils;

    function bit confirm(bit val);
        return val;
    endfunction

endpackage
