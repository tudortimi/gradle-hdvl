package main;
  import utils::*;
endpackage
