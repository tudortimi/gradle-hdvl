package some_published_dependency;
    `include "some_class.svh"
endpackage
