package uvc0;
endpackage
