package dummy;
endpackage
