module some_unit_test;
endmodule
