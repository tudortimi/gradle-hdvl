package some_package;

  `include "some_class.svh"

endpackage
