package some_other_package;

  `include "some_class.svh"

endpackage
