package proj1;
    import proj0::*;
endpackage
