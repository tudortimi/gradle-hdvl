class some_class;
endclass
