`define some_published_dependency_macro \
    $display("Hello from macro");
